* C:\Users\aryas\eSim-Workspace\switch_A\Counter_JK_3Nov.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 11/07/24 18:44:40

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  LOGIC_1 LOGIC_1 CLOCK Net-_U10-Pad4_ Net-_U10-Pad5_ Net-_U10-Pad3_ Net-_U5-Pad7_ d_jkff		
U10  Net-_U10-Pad1_ Net-_U10-Pad1_ Net-_U10-Pad3_ Net-_U10-Pad4_ Net-_U10-Pad5_ Net-_U10-Pad6_ Net-_U10-Pad7_ d_jkff		
v1  Net-_U1-Pad1_ GND pulse		
U1  Net-_U1-Pad1_ CLOCK adc_bridge_1		
v2  Net-_U3-Pad1_ GND DC		
U3  Net-_U3-Pad1_ LOGIC_1 adc_bridge_1		
U7  Net-_U10-Pad3_ Q0 dac_bridge_1		
U6  Net-_U5-Pad7_ Q0_bar dac_bridge_1		
U11  Net-_U10-Pad6_ Q1 dac_bridge_1		
U12  Net-_U10-Pad7_ Net-_R3-Pad1_ dac_bridge_1		
R2  Q0 GND 1k		
R4  Q1 GND 1k		
R1  Q0_bar GND 1k		
R3  Net-_R3-Pad1_ GND 1k		
U2  CLOCK plot_v1		
U4  LOGIC_1 plot_v1		
U9  Q0 plot_v1		
U8  Q0_bar plot_v1		
U14  Q1 plot_v1		
U13  Q1_bar plot_v1		
v3  Net-_U15-Pad1_ GND DC		
U15  Net-_U15-Pad1_ Net-_U10-Pad1_ adc_bridge_1		
U16  Net-_U10-Pad3_ Net-_U10-Pad6_ Net-_U16-Pad3_ d_xor		
U17  Net-_U16-Pad3_ Gray0 dac_bridge_1		
R5  Gray0 GND 1k		
U18  Gray0 plot_v1		

.end
